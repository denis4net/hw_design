library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity MEMCELL is
begin
	A, I, NRCK: in std_logic;
	O: out std_logic;
end MEMCELL;